`define STATE_RESET 3'h0
`define STATE_IF    3'h1
`define STATE_ID    3'h2
`define STATE_EX    3'h3