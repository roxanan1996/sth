`define OPSEL_NONE  3'h0
`define OPSEL_AND   3'h1
`define OPSEL_OR    3'h2
`define OPSEL_XOR   3'h3
`define OPSEL_NEG   3'h4
`define OPSEL_ADD   3'h5
`define OPSEL_SUB   3'h6
`define OPSEL_MUL   3'h7