module adder_subtractor(
    output  [3:0]   R,
    input   [3:0]   A,
    input   [3:0]   B,
    input           button
    );

    // TODO
endmodule
