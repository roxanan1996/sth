`define INSTRUCTION_NOP 16'h0000
`define INSTRUCTION_AND 16'h0001
`define INSTRUCTION_OR  16'h0002
`define INSTRUCTION_XOR 16'h0003
`define INSTRUCTION_NEG 16'h0004
`define INSTRUCTION_ADD 16'h0005
`define INSTRUCTION_SUB 16'h0006
`define INSTRUCTION_MUL 16'h0007